/*
The section of the CPU containing the register file, data memory, and ALU.
*/

module core (

);

// code here

endmodule