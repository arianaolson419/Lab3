/*
The section of the CPU containing the register file, data memory, and ALU.
*/

module core (
	input clk,
	input [31:0] rd,
	input [31:0] rt,
	input [31:0] rs,
	input [15:0] immediate,
	input [31:0] added_PC,
	output [31:0] Da,
	output is_zero
);

// code here

endmodule